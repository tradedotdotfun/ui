<svg width="24" height="24" viewBox="0 0 24 24" fill="currentColor" xmlns="http://www.w3.org/2000/svg">
<path d="M22 9.5L22 4.5L2 4.5L2 9.5L4.85714 9.5L4.85714 14.5L7.71428 14.5L7.71428 17L10.5714 17L10.5714 19.5L13.4286 19.5L13.4286 17L16.2857 17L16.2857 14.5L19.1429 14.5L19.1429 9.5L22 9.5Z" fill="currentColor"/>
</svg>
